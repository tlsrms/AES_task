`timescale 1ns / 1ps

module SubBytes(
    input wire [127:0] data_in,    // 128-bit input state
    output wire [127:0] data_out  // 128-bit output state
);

    // Instantiate 16 Sbox modules for parallel processing
    Sbox sbox0 (.data_in(data_in[127:120]), .data_out(data_out[127:120]));
    Sbox sbox1 (.data_in(data_in[119:112]), .data_out(data_out[119:112]));
    Sbox sbox2 (.data_in(data_in[111:104]), .data_out(data_out[111:104]));
    Sbox sbox3 (.data_in(data_in[103:96]),  .data_out(data_out[103:96]));
    Sbox sbox4 (.data_in(data_in[95:88]),   .data_out(data_out[95:88]));
    Sbox sbox5 (.data_in(data_in[87:80]),   .data_out(data_out[87:80]));
    Sbox sbox6 (.data_in(data_in[79:72]),   .data_out(data_out[79:72]));
    Sbox sbox7 (.data_in(data_in[71:64]),   .data_out(data_out[71:64]));
    Sbox sbox8 (.data_in(data_in[63:56]),   .data_out(data_out[63:56]));
    Sbox sbox9 (.data_in(data_in[55:48]),   .data_out(data_out[55:48]));
    Sbox sbox10 (.data_in(data_in[47:40]),  .data_out(data_out[47:40]));
    Sbox sbox11 (.data_in(data_in[39:32]),  .data_out(data_out[39:32]));
    Sbox sbox12 (.data_in(data_in[31:24]),  .data_out(data_out[31:24]));
    Sbox sbox13 (.data_in(data_in[23:16]),  .data_out(data_out[23:16]));
    Sbox sbox14 (.data_in(data_in[15:8]),   .data_out(data_out[15:8]));
    Sbox sbox15 (.data_in(data_in[7:0]),    .data_out(data_out[7:0]));

endmodule